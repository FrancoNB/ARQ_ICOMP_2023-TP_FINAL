`ifndef __IF_ID_VH__
`define __IF_ID_VH__
    `include "if.vh"
    `include "id.vh"

    `define DEFAULT_INSTRUCTION_SIZE `ARQUITECTURE_BITS
`endif // __IF_ID_VH__