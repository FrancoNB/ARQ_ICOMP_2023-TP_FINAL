`ifndef __DEBUGGER_VH__
`define __DEBUGGER_VH__
    `include "common.vh"

    `define DEFAULT_DEBUGGER_UART_BUS_SIZE          8
    `define DEFAULT_DEBUGGER_REGISTER_SIZE          `ARQUITECTURE_BITS
    `define DEFAULT_DEBUGGER_MEMORY_SLOT_SIZE       `ARQUITECTURE_BITS
    `define DEFAULT_DEBUGGER_REGISTER_BANK_BUS_SIZE `DEFAULT_DEBUGGER_REGISTER_SIZE * 32
    `define DEFAULT_DEBUGGER_MEMORY_DATA_BUS_SIZE   `ARQUITECTURE_BITS * 64

    `define DEBUGGER_STATE_IDLE              4'b0000
    `define DEBUGGER_STATE_LOAD              4'b0001
    `define DEBUGGER_STATE_RUN               4'b0010
    `define DEBUGGER_STATE_PRINT_REGISTERS   4'b0011
    `define DEBUGGER_STATE_PRINT_MEMORY_DATA 4'b0100
    `define DEBUGGER_STATE_UART_WR           4'b0101
    `define DEBUGGER_STATE_UART_WR_RESET     4'b0110
    `define DEBUGGER_STATE_UART_RD           4'b0111
    `define DEBUGGER_STATE_UART_RD_RESET     4'b1000


    `define DEBUGGER_NO_CICLE_MASK                  8'b00000000
    `define DEBUGGER_NO_ADDRESS_MASK                8'b00000000

    `define DEBUGGER_ERROR_PREFIX                   8'b11111111
    `define DEBUGGER_INFO_PREFIX                    8'b00000000

    `define DEBUGGER_INFO_END_PROGRAM               32'b00000000000000000000000000000001

    `define DEBUGGER_ERROR_INSTRUCTION_MEMORY_FULL  32'b00000000000000000000000000000001
    `define DEBUGGER_ERROR_NO_PROGRAM_LOAD          32'b00000000000000000000000000000010
    `define DEBUGGER_ERROR_BAD_REGISTER_ADDRESS     32'b00000000000000000000000000000011
    `define DEBUGGER_ERROR_BAD_MEMORY_ADDRESS       32'b00000000000000000000000000000100
    `define DEBUGGER_ERROR_UNKNOWN_COMMAND          32'b00000000000000000000000000000101
    `define DEBUGGER_ERROR_ALREADY_PROGRAM_LOAD     32'b00000000000000000000000000000110

`endif // __DEBUGGER_VH__