`ifndef __REGISTER_PRINTER_VH__
`define __REGISTER_PRINTER_VH__
    `include "common.vh"

    `define DEFAULT_REGISTER_PRINTER_UART_BUS_SIZE          8
    `define DEFAULT_REGISTER_PRINTER_OUT_BUS_SIZE           `DEFAULT_REGISTER_PRINTER_UART_BUS_SIZE * 7
    `define DEFAULT_REGISTER_PRINTER_REGISTER_SIZE          `ARQUITECTURE_BITS
    `define DEFAULT_REGISTER_PRINTER_REGISTER_BANK_BUS_SIZE `DEFAULT_REGISTER_PRINTER_REGISTER_SIZE * 32

    `define REGISTER_PRINTER_STATE_IDLE    2'b00
    `define REGISTER_PRINTER_STATE_PRINT   2'b01
    `define REGISTER_PRINTER_STATE_WAIT_WR 2'b10

`endif // __REGISTER_PRINTER_VH__