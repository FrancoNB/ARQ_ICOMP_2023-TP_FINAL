`ifndef __UART_VH__
`define __UART_VH__
    `define DATA_BITS 8
    `define SB_TICKS  16
    `define DVSR_BIT  9
    `define DVSR      326
    `define FIFO_SIZE 8
`endif // __UART_VH__