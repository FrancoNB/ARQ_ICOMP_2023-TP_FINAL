`ifndef __INSTRUCTION_MEMORY_VH__
`define __INSTRUCTION_MEMORY_VH__
    `include "common.vh"

    `define DEFAULT_INSTRUCTION_MEMORY_REG_SIZE `ARQUITECTURE_BITS
    `define DEFAULT_INSTRUCTION_MEMORY_MEM_SIZE 320
    
    `define NUMBER_OF_STATE_INSTRUCTION_MEMORY        5
    `define BITS_FOR_STATE_COUNTER_INSTRUCTION_MEMORY $clog2(`NUMBER_OF_STATE_INSTRUCTION_MEMORY)

    `define STATE_INSTRUCTION_MEMORY_IDLE              3'b000
    `define STATE_INSTRUCTION_MEMORY_WRITE_INSTRUCTION 3'b001
    `define STATE_INSTRUCTION_MEMORY_READY_TO_EXECUTE  3'b010
    `define STATE_INSTRUCTION_MEMORY_SEND_INSTRUCTION  3'b011
    `define STATE_INSTRUCTION_PROGRAM_FINISHED         3'b100
`endif // __INSTRUCTION_MEMORY_VH__