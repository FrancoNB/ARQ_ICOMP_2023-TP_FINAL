`ifndef __INSTRUCTION_MEMORY_VH__
`define __INSTRUCTION_MEMORY_VH__
    `include "common.vh"

    `define DEFAULT_INSTRUCTION_MEMORY_WORD_SIZE_IN_BYTES `ARQUITECTURE_BITS / `BYTE_SIZE 
    `define DEFAULT_INSTRUCTION_MEMORY_MEM_SIZE_IN_WORDS  10
    
    `define NUMBER_OF_STATE_INSTRUCTION_MEMORY        2
    `define BITS_FOR_STATE_COUNTER_INSTRUCTION_MEMORY $clog2(`NUMBER_OF_STATE_INSTRUCTION_MEMORY)

    `define STATE_INSTRUCTION_MEMORY_WRITE 2'b0
    `define STATE_INSTRUCTION_MEMORY_READ  2'b1
`endif // __INSTRUCTION_MEMORY_VH__