`ifndef __TOP_VH__
`define __TOP_VH__
    `include "common.vh"
    `include "mips.vh"
    `include "debugger.vh"
    `include "uart.vh"
`endif // __TOP_VH__