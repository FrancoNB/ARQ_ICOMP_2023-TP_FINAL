`ifndef __ADDER_VH__
`define __ADDER_VH__
    `define DEFAULT_ADDER_BUS_SIZE 32
`endif // __ADDER_VH__