`ifndef __AND_VH__
`define __AND_VH__
    `include "common.vh"

    `define DEFAULT_AND_CHANNELS 2
`endif // __AND_VH__