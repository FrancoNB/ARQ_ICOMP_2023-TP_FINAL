`ifndef __MUX_VH__
`define __MUX_VH__
    `define DEFAULT_MUX_CHANNELS 2
    `define DEFAULT_MUX_BUS_SIZE 32
`endif // __MUX_VH__s